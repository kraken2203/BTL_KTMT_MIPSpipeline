library verilog;
use verilog.vl_types.all;
entity ALUDec_tb is
end ALUDec_tb;
