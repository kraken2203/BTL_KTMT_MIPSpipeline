library verilog;
use verilog.vl_types.all;
entity MainDec_tb is
end MainDec_tb;
