`timescale 10ns/1ns 
module RegFile_tb();
